
--******************************************************--
--        PONTIFICIA UNIVERSIDAD JAVERIANA              --
--                Disegno Digital                       --
--              PROYECTO CAJA FUERTE                    --
-- 							                            --
-- Titulo :    Sumador Decimal digito		            --
-- Fecha  :  	D:01 M:10 Y:2019                        --
--******************************************************--
